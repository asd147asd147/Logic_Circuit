module tFF_tb;

wire Q;
reg T;
reg clock;
reg reset;

tFF
 U0 (
  .Q(Q),
  .T(T),
  .clock(clock),
  .reset(reset));

  initial
  begin
    T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
    #100 T = 1'b0;
    #100 T = 1'b1;
  end

  initial
  begin
    clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
    #100 clock = 1'b0;
    #100 clock = 1'b1;
  end

  initial
  begin
    reset = 1'b1;
    #100 reset = 1'b0;
  end

endmodule
