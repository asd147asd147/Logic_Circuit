/***********************
*
* Jong-gyu Park
* pjk5401@gmail.com
* 2016/09/02
*
***********************/

module PNU_OR8(i1, i2, i3, i4, i5, i6, i7, i8, o1);
    input i1, i2, i3, i4, i5, i6, i7, i8;
    output o1;
    assign o1 = i1 | i2 | i3 | i4 | i5 | i6 | i7 | i8;
endmodule