/***********************
*
* Jong-gyu Park
* pjk5401@gmail.com
* 2016/09/02
*
***********************/

module PNU_ONE(o1);
    output o1;
    assign o1=1;
endmodule